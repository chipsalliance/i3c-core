// SPDX-License-Identifier: Apache-2.0

// Command Queue for I3C Controller Interface
module cmd_queue #() (
    // TODO: Provide Command Queue Interface
    // see https://github.com/lowRISC/opentitan/blob/c97dc79d6fef6b30929a0b7da9e2c4dbc653711c/hw/ip/i2c/rtl/i2c_controller_fsm.sv#L22
    // for reference
);
endmodule
