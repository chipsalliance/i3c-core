`include "base_vseq.sv"
`include "direct_vseq.sv"
`include "direct_with_rstart_vseq.sv"
`include "broadcast_followed_by_data_vseq.sv"
`include "broadcast_followed_by_data_with_rstart_vseq.sv"
`include "direct_i2c_vseq.sv"
`include "direct_i2c_with_rstart_vseq.sv"
`include "broadcast_followed_by_i2c_data_vseq.sv"
`include "broadcast_followed_by_i2c_data_with_rstart_vseq.sv"
