package i3c_sequence_env_pkg;
  import uvm_pkg::*;
  import i3c_agent_pkg::*;


  `include "i3c_sequence_env_cfg.sv"
  `include "i3c_sequence_env.sv"
endpackage
