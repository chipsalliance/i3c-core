package i3c_sequence_env_pkg;
  import uvm_pkg::*;
  import i3c_agent_pkg::*;

  typedef class i3c_sequence_virtual_sequencer;
  `include "i3c_sequence_env_cfg.sv"
  `include "i3c_sequence_virtual_sequencer.sv"
  `include "i3c_sequence_env.sv"
  `include "i3c_base_vseq.sv"
  `include "i3c_sequence_vseq_list.sv"
endpackage
