// Copyright (c) 2024 Antmicro <www.antmicro.com>
// SPDX-License-Identifier: Apache-2.0

package i3c_ctrl_pkg;

  // To raise errors
  typedef struct packed {logic err_0;} i3c_err_t;

  // To raise interrupts
  typedef struct packed {logic irq_0;} i3c_irq_t;

  // I3C Packet
  typedef struct packed {logic irq_0;} i3c_ah_t;

endpackage
