package i3c_sequence_test_pkg;
  import uvm_pkg::*;
  import i3c_sequence_env_pkg::*;

  `include "i3c_sequence_test.sv"
endpackage
