`include "i3c_sequence_direct_vseq.sv"
