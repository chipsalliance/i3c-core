package i3c_test_pkg;
  // dep packages
  import uvm_pkg::*;
  import i3c_env_pkg::*;

  `include "i3c_base_test.sv"

endpackage

