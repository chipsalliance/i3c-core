`include "i3c_base_vseq.sv"
