`include "i3c_direct_data_seq.sv"
`include "i3c_direct_data_with_rstart_seq.sv"
`include "i3c_broadcast_followed_by_data_seq.sv"
`include "i3c_broadcast_followed_by_data_with_rstart_seq.sv"
`include "i2c_direct_data_seq.sv"
`include "i2c_direct_data_with_rstart_seq.sv"
`include "i3c_broadcast_followed_by_i2c_data_seq.sv"
`include "i3c_broadcast_followed_by_i2c_data_with_rstart_seq.sv"
