package i3c_test_pkg;
  // dep packages
  import uvm_pkg::*;
  import i3c_env_pkg::*;

  `include "uvm_macros.svh"

  `include "i3c_base_test.sv"

endpackage

