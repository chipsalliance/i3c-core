`include "i3c_direct_data_seq.sv"
`include "i3c_direct_data_with_repeated_start_seq.sv"
`include "i3c_broadcast_followed_by_data_seq.sv"
