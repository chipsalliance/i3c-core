`include "i3c_base_seq.sv"
