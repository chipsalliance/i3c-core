`include "i3c_sequence_base_vseq.sv"
`include "i3c_sequence_direct_vseq.sv"
`include "i3c_sequence_direct_with_repeated_start_vseq.sv"
